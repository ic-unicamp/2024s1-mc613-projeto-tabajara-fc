module movimento (
    input reset,
    input btn_D,
    output posX,

)