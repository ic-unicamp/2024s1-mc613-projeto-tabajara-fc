module tela_inicial(
    input reset,
    input [9:0] h_counter,
    input [9:0] v_counter,
    output reg [7:0] R,
    output reg [7:8] G,
    output reg [7:8] B
);


endmodule